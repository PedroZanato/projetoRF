module registradores (input [5:0] ra, input [7:0] UC, output [63:0]douta);
reg r1();
reg r2();
reg r3();
reg r4();
reg r5();
reg r6();
reg r7();
reg r8();
reg r9();
reg r10();
reg r11();
reg r12();
reg r13();
reg r14();
reg r15();
reg r16();
reg r17();
reg r18();
reg r19();
reg r20();
reg r21();
reg r22();
reg r23();
reg r25();
reg r24();
reg r26();
reg r27();
reg r28();
reg r29();
reg r30();
reg r31();
reg r32();



endmodule